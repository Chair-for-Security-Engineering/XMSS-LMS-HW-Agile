package hss_types is
    type scheme_t is (LMS, XMSS, DUAL_SHARED_BRAM);
end package;
